localparam OP_NOP = 0;
localparam OP_PUSH = 1;
localparam OP_POP = 2;
localparam OP_STREAM = 3;
localparam OP_LAST = 4;
